module control_unit(instruction, status, reset, clock, controlWord, K);
    parameter cw_bits = 31;
    parameter K_bits = 64;
    input [31:0] instruction;
    input [4:0] status;     // V, C, N, Z
    input reset, clock;
    output [cw_bits-1:0] controlWord;
    output [K_bits-1:0] K;
    
    wire [10:0] opcode;
    
    assign opcode = instruction[31:21];
    
    // partial control words
    wire [cw_bits+K_bits+1:0] branch_cw, other_cw;
    
    // controlWord
    wire [cw_bits-1:0] D_Transfer_cw, I_Arithmetic_cw, I_Logic_cw, IW_cw, R_ALU_cw;
    wire [cw_bits-1:0] B_cw, B_conditional_cw, BL_cw, CBZ_CBNZ_cw, BR_cw;
    
    // nextState
    wire [1:0] D_Transfer_ns, I_Arithmetic_ns, I_Logic_ns, IW_ns, R_ALU_ns;
    wire [1:0] B_ns, B_conditional_ns, BL_ns, CBZ_CBNZ_ns, BR_ns;
    
    // K
    wire [K_bits-1:0] D_Transfer_K, I_Arithmetic_K, I_Logic_K, IW_K, R_ALU_K;
    wire [K_bits-1:0] B_K, B_conditional_K, BL_K, CBZ_CBNZ_K, BR_K;
    
    // concatenated controlWord + K + nextState
    wire [cw_bits+K_bits+1:0] D_Transfer_cwc, I_Arithmetic_cwc, I_Logic_cwc, IW_cwc, R_ALU_cwc;
    wire [cw_bits+K_bits+1:0] B_cwc, B_conditional_cwc, BL_cwc, CBZ_CBNZ_cwc, BR_cwc;
    
    // state logic
    wire [1:0] nextState;
    reg [1:0] state;
    always @(posedge clock or posedge reset) begin
        if(reset)
            state <= 2'b00;
        else
            state <= nextState;
    end
    
    // decoder module definitions
    B dec1_000 (instruction, state, B_cw, B_ns, B_K);
    assign B_cwc = {B_cw, B_K, B_ns};
    B_cond dec1_010 (status, instruction, state, B_conditional_cw, B_conditional_ns, B_conditional_K);
    assign B_conditional_cwc = {B_conditional_cw, B_conditional_K, B_conditional_ns};
    B_link dec1_100 (instruction, state, BL_cw, BL_ns, BL_K);
    assign BL_cwc = {BL_cw, BL_K, BL_ns};
    B_compare dec1_101 (status, instruction, state, CBZ_CBNZ_cw, CBZ_CBNZ_ns, CBZ_CBNZ_K);
    assign CBZ_CBNZ_cwc = {CBZ_CBNZ_cw, CBZ_CBNZ_K, CBZ_CBNZ_ns};
    B_to_reg dec1_110 (instruction, state, BR_cw, BR_ns, BR_K);
    assign BR_cwc = {BR_cw, BR_K, BR_ns};
    
    D dec0_000 (instruction, state, D_Transfer_cw, D_Transfer_ns, D_Transfer_K);
    assign D_Transfer_cwc = {D_Transfer_cw, D_Transfer_K, D_Transfer_ns};
    I_arithmetic dec0_010 (instruction, state, I_Arithmetic_cw, I_Arithmetic_ns, I_Arithmetic_K);
    assign I_Arithmetic_cwc = {I_Arithmetic_cw, I_Arithmetic_K, I_Arithmetic_ns};
    I_logic dec0_100 (instruction, state, I_Logic_cw, I_Logic_ns, I_Logic_K);
    assign I_Logic_cwc = {I_Logic_cw, I_Logic_K, I_Logic_ns};
    WI dec0_101 (instruction, state, IW_cw, IW_ns, IW_K);
    assign IW_cwc = {IW_cw, IW_K, IW_ns};
    R dec0_110 (instruction, state, R_ALU_cw, R_ALU_ns, R_ALU_K);
    assign R_ALU_cwc = {R_ALU_cw, R_ALU_K, R_ALU_ns};
    
    // 8:1 mux to select between branch instructions
    Mux8to1Nbit branch_mux (opcode[10:8],
        B_cwc, 0, B_conditional_cwc, 0, BL_cwc,
        CBZ_CBNZ_cwc, BR_cwc, 0, branch_cw);
    defparam branch_mux.N = (cw_bits+K_bits+2);
    
    // 8:1 mux to select between all other instructions
    Mux8to1Nbit other_mux (opcode[4:2],
        D_Transfer_cwc, 0, I_Arithmetic_cwc, 0, I_Logic_cwc,
        IW_cwc, R_ALU_cwc, 0, other_cw);
    defparam other_mux.N = (cw_bits+K_bits+2);
    
    // 2:1 mux to select between branch instructions and all others
    assign controlWord = opcode[5] ? branch_cw[cw_bits+K_bits+1:K_bits+2] : other_cw[cw_bits+K_bits+1:K_bits+2];
    assign K = opcode[5] ? branch_cw[K_bits+1:2] : other_cw[K_bits+1:2];
    assign nextState = opcode[5] ? branch_cw[1:0] : other_cw[1:0];
    
endmodule